
# Created      : Thu May 23 15:40:21 2002
# Platform     : Linux 2.4.10 #1 Fri Sep 28 09:29:45 EDT 2001 i686 
# User         : sadya@voskhod.eecs.umich.edu (Saurabh N Adya,Not Available,NotAvailable/Freysinger;CR0i;30) 

NAMESCASESENSITIVE ON ;
UNITS
DATABASE MICRONS 100 ;
END UNITS

LAYER poly
	TYPE MASTERSLICE ;
END poly
LAYER cont
	TYPE CUT ;
END cont
LAYER metal1
	TYPE ROUTING ;
	PITCH 1.7 ;
	WIDTH .8 ;
	SPACING .6 ;
	DIRECTION HORIZONTAL ;
END metal1

LAYER via1
	TYPE CUT ;
END via1

LAYER metal2
	TYPE ROUTING ;
	PITCH 2 ;
	WIDTH .8 ;
	SPACING .9 ;
	DIRECTION VERTICAL ;
END metal2

LAYER via2
	TYPE CUT ;
END via2

LAYER metal3
	TYPE ROUTING ;
	PITCH 1.7 ;
	WIDTH .8 ;
	SPACING .9 ;
	DIRECTION HORIZONTAL ;
END metal3

LAYER OVERLAP
	TYPE OVERLAP ;
END OVERLAP
VIA cont DEFAULT
	LAYER poly ;
		RECT -.6 -.6 .6 .6 ;
	LAYER cont ;
		RECT -.3 -.3 .3 .3 ;
	LAYER metal1 ;
		RECT -.4 -.4 .4 .4 ;
END cont

VIA via1 DEFAULT
	LAYER metal1 ;
		RECT -.7 -.7 .7 .7 ;
	LAYER via1 ;
		RECT -.3 -.3 .3 .3 ;
	LAYER metal2 ;
		RECT -.4 -.4 .4 .4 ;
END via1

VIA via2 DEFAULT
	LAYER metal2 ;
		RECT -.65 -.65 .65 .65 ;
	LAYER via2 ;
		RECT -.3 -.3 .3 .3 ;
	LAYER metal3 ;
		RECT -.4 -.4 .4 .4 ;
END via2

SPACING
	SAMENET metal1 metal1 .6 ;
	SAMENET metal2 metal2 .9 ;
	SAMENET metal3 metal3 .9 ;
	SAMENET cont cont .8 ;
	SAMENET cont via1 .65 ;
	SAMENET via1 via1 1 ;
	SAMENET via1 via2 .6 ;
	SAMENET via2 via1 1 ;
END SPACING
SITE core
	SIZE 0.01 BY 0.16 ;
	CLASS CORE ;
	SYMMETRY  Y  ;
END core

MACRO MAS0
	CLASS CORE ;
	SIZE 0.01 BY 0.01 ;
	ORIGIN 0 0 ;
	SYMMETRY X ;
	SITE core 0 0 N DO 1 BY 1 STEP 0 0 ;
	PIN P1
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.00495 0.00495 0.00505 0.00505 ;
		END
	END P1
END MAS0

MACRO MAS1
	CLASS CORE ;
	SIZE 0.02 BY 0.16 ;
	ORIGIN 0 0 ;
	SYMMETRY X ;
	SITE core 0 0 N DO 1 BY 1 STEP 0 0 ;
	PIN P1
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0099 0.0792 0.0101 0.0808 ;
		END
	END P1
END MAS1

MACRO MAS2
	CLASS CORE ;
	SIZE 0.02 BY 0.16 ;
	ORIGIN 0 0 ;
	SYMMETRY X ;
	SITE core 0 0 N DO 1 BY 1 STEP 0 0 ;
	PIN P1
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0099 0.0792 0.0101 0.0808 ;
		END
	END P1
	PIN P2
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0099 0.0792 0.0101 0.0808 ;
		END
	END P2
END MAS2

MACRO MAS3
	CLASS CORE ;
	SIZE 0.04 BY 0.16 ;
	ORIGIN 0 0 ;
	SYMMETRY X ;
	SITE core 0 0 N DO 1 BY 1 STEP 0 0 ;
	PIN P1
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0198 0.0792 0.0202 0.0808 ;
		END
	END P1
END MAS3

MACRO MAS4
	CLASS CORE ;
	SIZE 0.04 BY 0.16 ;
	ORIGIN 0 0 ;
	SYMMETRY X ;
	SITE core 0 0 N DO 1 BY 1 STEP 0 0 ;
	PIN P1
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0198 0.0792 0.0202 0.0808 ;
		END
	END P1
	PIN P2
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0198 0.0792 0.0202 0.0808 ;
		END
	END P2
END MAS4

MACRO MAS5
	CLASS CORE ;
	SIZE 0.04 BY 0.16 ;
	ORIGIN 0 0 ;
	SYMMETRY X ;
	SITE core 0 0 N DO 1 BY 1 STEP 0 0 ;
	PIN P1
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0198 0.0792 0.0202 0.0808 ;
		END
	END P1
	PIN P2
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0198 0.0792 0.0202 0.0808 ;
		END
	END P2
	PIN P3
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0198 0.0792 0.0202 0.0808 ;
		END
	END P3
END MAS5

MACRO MAS6
	CLASS CORE ;
	SIZE 0.06 BY 0.16 ;
	ORIGIN 0 0 ;
	SYMMETRY X ;
	SITE core 0 0 N DO 1 BY 1 STEP 0 0 ;
	PIN P1
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0297 0.0792 0.0303 0.0808 ;
		END
	END P1
	PIN P2
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0297 0.0792 0.0303 0.0808 ;
		END
	END P2
END MAS6

MACRO MAS7
	CLASS CORE ;
	SIZE 0.06 BY 0.16 ;
	ORIGIN 0 0 ;
	SYMMETRY X ;
	SITE core 0 0 N DO 1 BY 1 STEP 0 0 ;
	PIN P1
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0297 0.0792 0.0303 0.0808 ;
		END
	END P1
	PIN P2
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0297 0.0792 0.0303 0.0808 ;
		END
	END P2
	PIN P3
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0297 0.0792 0.0303 0.0808 ;
		END
	END P3
END MAS7

MACRO MAS8
	CLASS CORE ;
	SIZE 0.06 BY 0.16 ;
	ORIGIN 0 0 ;
	SYMMETRY X ;
	SITE core 0 0 N DO 1 BY 1 STEP 0 0 ;
	PIN P1
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0297 0.0792 0.0303 0.0808 ;
		END
	END P1
	PIN P2
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0297 0.0792 0.0303 0.0808 ;
		END
	END P2
	PIN P3
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0297 0.0792 0.0303 0.0808 ;
		END
	END P3
	PIN P4
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0297 0.0792 0.0303 0.0808 ;
		END
	END P4
END MAS8

MACRO MAS9
	CLASS CORE ;
	SIZE 0.06 BY 0.16 ;
	ORIGIN 0 0 ;
	SYMMETRY X ;
	SITE core 0 0 N DO 1 BY 1 STEP 0 0 ;
	PIN P1
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0297 0.0792 0.0303 0.0808 ;
		END
	END P1
	PIN P2
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0297 0.0792 0.0303 0.0808 ;
		END
	END P2
	PIN P3
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0297 0.0792 0.0303 0.0808 ;
		END
	END P3
	PIN P4
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0297 0.0792 0.0303 0.0808 ;
		END
	END P4
	PIN P5
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0297 0.0792 0.0303 0.0808 ;
		END
	END P5
END MAS9

MACRO MAS10
	CLASS CORE ;
	SIZE 0.08 BY 0.16 ;
	ORIGIN 0 0 ;
	SYMMETRY X ;
	SITE core 0 0 N DO 1 BY 1 STEP 0 0 ;
	PIN P1
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0396 0.0792 0.0404 0.0808 ;
		END
	END P1
END MAS10

MACRO MAS11
	CLASS CORE ;
	SIZE 0.08 BY 0.16 ;
	ORIGIN 0 0 ;
	SYMMETRY X ;
	SITE core 0 0 N DO 1 BY 1 STEP 0 0 ;
	PIN P1
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0396 0.0792 0.0404 0.0808 ;
		END
	END P1
	PIN P2
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0396 0.0792 0.0404 0.0808 ;
		END
	END P2
END MAS11

MACRO MAS12
	CLASS CORE ;
	SIZE 0.08 BY 0.16 ;
	ORIGIN 0 0 ;
	SYMMETRY X ;
	SITE core 0 0 N DO 1 BY 1 STEP 0 0 ;
	PIN P1
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0396 0.0792 0.0404 0.0808 ;
		END
	END P1
	PIN P2
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0396 0.0792 0.0404 0.0808 ;
		END
	END P2
	PIN P3
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0396 0.0792 0.0404 0.0808 ;
		END
	END P3
END MAS12

MACRO MAS13
	CLASS CORE ;
	SIZE 0.08 BY 0.16 ;
	ORIGIN 0 0 ;
	SYMMETRY X ;
	SITE core 0 0 N DO 1 BY 1 STEP 0 0 ;
	PIN P1
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0396 0.0792 0.0404 0.0808 ;
		END
	END P1
	PIN P2
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0396 0.0792 0.0404 0.0808 ;
		END
	END P2
	PIN P3
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0396 0.0792 0.0404 0.0808 ;
		END
	END P3
	PIN P4
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0396 0.0792 0.0404 0.0808 ;
		END
	END P4
END MAS13

MACRO MAS14
	CLASS CORE ;
	SIZE 0.08 BY 0.16 ;
	ORIGIN 0 0 ;
	SYMMETRY X ;
	SITE core 0 0 N DO 1 BY 1 STEP 0 0 ;
	PIN P1
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0396 0.0792 0.0404 0.0808 ;
		END
	END P1
	PIN P2
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0396 0.0792 0.0404 0.0808 ;
		END
	END P2
	PIN P3
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0396 0.0792 0.0404 0.0808 ;
		END
	END P3
	PIN P4
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0396 0.0792 0.0404 0.0808 ;
		END
	END P4
	PIN P5
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0396 0.0792 0.0404 0.0808 ;
		END
	END P5
END MAS14

MACRO MAS15
	CLASS CORE ;
	SIZE 0.1 BY 0.16 ;
	ORIGIN 0 0 ;
	SYMMETRY X ;
	SITE core 0 0 N DO 1 BY 1 STEP 0 0 ;
	PIN P1
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0495 0.0792 0.0505 0.0808 ;
		END
	END P1
	PIN P2
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0495 0.0792 0.0505 0.0808 ;
		END
	END P2
END MAS15

MACRO MAS16
	CLASS CORE ;
	SIZE 0.1 BY 0.16 ;
	ORIGIN 0 0 ;
	SYMMETRY X ;
	SITE core 0 0 N DO 1 BY 1 STEP 0 0 ;
	PIN P1
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0495 0.0792 0.0505 0.0808 ;
		END
	END P1
	PIN P2
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0495 0.0792 0.0505 0.0808 ;
		END
	END P2
	PIN P3
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0495 0.0792 0.0505 0.0808 ;
		END
	END P3
	PIN P4
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0495 0.0792 0.0505 0.0808 ;
		END
	END P4
END MAS16

MACRO MAS17
	CLASS CORE ;
	SIZE 0.1 BY 0.16 ;
	ORIGIN 0 0 ;
	SYMMETRY X ;
	SITE core 0 0 N DO 1 BY 1 STEP 0 0 ;
	PIN P1
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0495 0.0792 0.0505 0.0808 ;
		END
	END P1
	PIN P2
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0495 0.0792 0.0505 0.0808 ;
		END
	END P2
	PIN P3
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0495 0.0792 0.0505 0.0808 ;
		END
	END P3
	PIN P4
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0495 0.0792 0.0505 0.0808 ;
		END
	END P4
	PIN P5
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0495 0.0792 0.0505 0.0808 ;
		END
	END P5
END MAS17

MACRO MAS18
	CLASS CORE ;
	SIZE 0.1 BY 0.16 ;
	ORIGIN 0 0 ;
	SYMMETRY X ;
	SITE core 0 0 N DO 1 BY 1 STEP 0 0 ;
	PIN P1
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0495 0.0792 0.0505 0.0808 ;
		END
	END P1
	PIN P2
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0495 0.0792 0.0505 0.0808 ;
		END
	END P2
	PIN P3
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0495 0.0792 0.0505 0.0808 ;
		END
	END P3
	PIN P4
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0495 0.0792 0.0505 0.0808 ;
		END
	END P4
	PIN P5
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0495 0.0792 0.0505 0.0808 ;
		END
	END P5
	PIN P6
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0495 0.0792 0.0505 0.0808 ;
		END
	END P6
END MAS18

MACRO MAS19
	CLASS CORE ;
	SIZE 0.1 BY 0.16 ;
	ORIGIN 0 0 ;
	SYMMETRY X ;
	SITE core 0 0 N DO 1 BY 1 STEP 0 0 ;
	PIN P1
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0495 0.0792 0.0505 0.0808 ;
		END
	END P1
	PIN P2
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0495 0.0792 0.0505 0.0808 ;
		END
	END P2
	PIN P3
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0495 0.0792 0.0505 0.0808 ;
		END
	END P3
	PIN P4
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0495 0.0792 0.0505 0.0808 ;
		END
	END P4
	PIN P5
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0495 0.0792 0.0505 0.0808 ;
		END
	END P5
	PIN P6
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0495 0.0792 0.0505 0.0808 ;
		END
	END P6
	PIN P7
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0495 0.0792 0.0505 0.0808 ;
		END
	END P7
END MAS19

MACRO MAS20
	CLASS CORE ;
	SIZE 0.12 BY 0.16 ;
	ORIGIN 0 0 ;
	SYMMETRY X ;
	SITE core 0 0 N DO 1 BY 1 STEP 0 0 ;
	PIN P1
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0594 0.0792 0.0606 0.0808 ;
		END
	END P1
	PIN P2
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0594 0.0792 0.0606 0.0808 ;
		END
	END P2
END MAS20

MACRO MAS21
	CLASS CORE ;
	SIZE 0.12 BY 0.16 ;
	ORIGIN 0 0 ;
	SYMMETRY X ;
	SITE core 0 0 N DO 1 BY 1 STEP 0 0 ;
	PIN P1
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0594 0.0792 0.0606 0.0808 ;
		END
	END P1
	PIN P2
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0594 0.0792 0.0606 0.0808 ;
		END
	END P2
	PIN P3
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0594 0.0792 0.0606 0.0808 ;
		END
	END P3
END MAS21

MACRO MAS22
	CLASS CORE ;
	SIZE 0.12 BY 0.16 ;
	ORIGIN 0 0 ;
	SYMMETRY X ;
	SITE core 0 0 N DO 1 BY 1 STEP 0 0 ;
	PIN P1
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0594 0.0792 0.0606 0.0808 ;
		END
	END P1
	PIN P2
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0594 0.0792 0.0606 0.0808 ;
		END
	END P2
	PIN P3
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0594 0.0792 0.0606 0.0808 ;
		END
	END P3
	PIN P4
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0594 0.0792 0.0606 0.0808 ;
		END
	END P4
END MAS22

MACRO MAS23
	CLASS CORE ;
	SIZE 0.12 BY 0.16 ;
	ORIGIN 0 0 ;
	SYMMETRY X ;
	SITE core 0 0 N DO 1 BY 1 STEP 0 0 ;
	PIN P1
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0594 0.0792 0.0606 0.0808 ;
		END
	END P1
	PIN P2
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0594 0.0792 0.0606 0.0808 ;
		END
	END P2
	PIN P3
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0594 0.0792 0.0606 0.0808 ;
		END
	END P3
	PIN P4
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0594 0.0792 0.0606 0.0808 ;
		END
	END P4
	PIN P5
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0594 0.0792 0.0606 0.0808 ;
		END
	END P5
END MAS23

MACRO MAS24
	CLASS CORE ;
	SIZE 0.12 BY 0.16 ;
	ORIGIN 0 0 ;
	SYMMETRY X ;
	SITE core 0 0 N DO 1 BY 1 STEP 0 0 ;
	PIN P1
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0594 0.0792 0.0606 0.0808 ;
		END
	END P1
	PIN P2
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0594 0.0792 0.0606 0.0808 ;
		END
	END P2
	PIN P3
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0594 0.0792 0.0606 0.0808 ;
		END
	END P3
	PIN P4
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0594 0.0792 0.0606 0.0808 ;
		END
	END P4
	PIN P5
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0594 0.0792 0.0606 0.0808 ;
		END
	END P5
	PIN P6
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0594 0.0792 0.0606 0.0808 ;
		END
	END P6
END MAS24

MACRO MAS25
	CLASS CORE ;
	SIZE 0.12 BY 0.16 ;
	ORIGIN 0 0 ;
	SYMMETRY X ;
	SITE core 0 0 N DO 1 BY 1 STEP 0 0 ;
	PIN P1
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0594 0.0792 0.0606 0.0808 ;
		END
	END P1
	PIN P2
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0594 0.0792 0.0606 0.0808 ;
		END
	END P2
	PIN P3
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0594 0.0792 0.0606 0.0808 ;
		END
	END P3
	PIN P4
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0594 0.0792 0.0606 0.0808 ;
		END
	END P4
	PIN P5
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0594 0.0792 0.0606 0.0808 ;
		END
	END P5
	PIN P6
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0594 0.0792 0.0606 0.0808 ;
		END
	END P6
	PIN P7
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0594 0.0792 0.0606 0.0808 ;
		END
	END P7
END MAS25

MACRO MAS26
	CLASS CORE ;
	SIZE 0.12 BY 0.16 ;
	ORIGIN 0 0 ;
	SYMMETRY X ;
	SITE core 0 0 N DO 1 BY 1 STEP 0 0 ;
	PIN P1
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0594 0.0792 0.0606 0.0808 ;
		END
	END P1
	PIN P2
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0594 0.0792 0.0606 0.0808 ;
		END
	END P2
	PIN P3
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0594 0.0792 0.0606 0.0808 ;
		END
	END P3
	PIN P4
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0594 0.0792 0.0606 0.0808 ;
		END
	END P4
	PIN P5
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0594 0.0792 0.0606 0.0808 ;
		END
	END P5
	PIN P6
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0594 0.0792 0.0606 0.0808 ;
		END
	END P6
	PIN P7
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0594 0.0792 0.0606 0.0808 ;
		END
	END P7
	PIN P8
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0594 0.0792 0.0606 0.0808 ;
		END
	END P8
END MAS26

MACRO MAS27
	CLASS CORE ;
	SIZE 0.12 BY 0.16 ;
	ORIGIN 0 0 ;
	SYMMETRY X ;
	SITE core 0 0 N DO 1 BY 1 STEP 0 0 ;
	PIN P1
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0594 0.0792 0.0606 0.0808 ;
		END
	END P1
	PIN P2
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0594 0.0792 0.0606 0.0808 ;
		END
	END P2
	PIN P3
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0594 0.0792 0.0606 0.0808 ;
		END
	END P3
	PIN P4
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0594 0.0792 0.0606 0.0808 ;
		END
	END P4
	PIN P5
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0594 0.0792 0.0606 0.0808 ;
		END
	END P5
	PIN P6
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0594 0.0792 0.0606 0.0808 ;
		END
	END P6
	PIN P7
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0594 0.0792 0.0606 0.0808 ;
		END
	END P7
	PIN P8
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0594 0.0792 0.0606 0.0808 ;
		END
	END P8
	PIN P9
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0594 0.0792 0.0606 0.0808 ;
		END
	END P9
END MAS27

MACRO MAS28
	CLASS CORE ;
	SIZE 0.14 BY 0.16 ;
	ORIGIN 0 0 ;
	SYMMETRY X ;
	SITE core 0 0 N DO 1 BY 1 STEP 0 0 ;
	PIN P1
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0693 0.0792 0.0707 0.0808 ;
		END
	END P1
	PIN P2
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0693 0.0792 0.0707 0.0808 ;
		END
	END P2
END MAS28

MACRO MAS29
	CLASS CORE ;
	SIZE 0.14 BY 0.16 ;
	ORIGIN 0 0 ;
	SYMMETRY X ;
	SITE core 0 0 N DO 1 BY 1 STEP 0 0 ;
	PIN P1
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0693 0.0792 0.0707 0.0808 ;
		END
	END P1
	PIN P2
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0693 0.0792 0.0707 0.0808 ;
		END
	END P2
	PIN P3
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0693 0.0792 0.0707 0.0808 ;
		END
	END P3
	PIN P4
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0693 0.0792 0.0707 0.0808 ;
		END
	END P4
END MAS29

MACRO MAS30
	CLASS CORE ;
	SIZE 0.14 BY 0.16 ;
	ORIGIN 0 0 ;
	SYMMETRY X ;
	SITE core 0 0 N DO 1 BY 1 STEP 0 0 ;
	PIN P1
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0693 0.0792 0.0707 0.0808 ;
		END
	END P1
	PIN P2
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0693 0.0792 0.0707 0.0808 ;
		END
	END P2
	PIN P3
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0693 0.0792 0.0707 0.0808 ;
		END
	END P3
	PIN P4
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0693 0.0792 0.0707 0.0808 ;
		END
	END P4
	PIN P5
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0693 0.0792 0.0707 0.0808 ;
		END
	END P5
END MAS30

MACRO MAS31
	CLASS CORE ;
	SIZE 0.14 BY 0.16 ;
	ORIGIN 0 0 ;
	SYMMETRY X ;
	SITE core 0 0 N DO 1 BY 1 STEP 0 0 ;
	PIN P1
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0693 0.0792 0.0707 0.0808 ;
		END
	END P1
	PIN P2
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0693 0.0792 0.0707 0.0808 ;
		END
	END P2
	PIN P3
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0693 0.0792 0.0707 0.0808 ;
		END
	END P3
	PIN P4
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0693 0.0792 0.0707 0.0808 ;
		END
	END P4
	PIN P5
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0693 0.0792 0.0707 0.0808 ;
		END
	END P5
	PIN P6
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0693 0.0792 0.0707 0.0808 ;
		END
	END P6
END MAS31

MACRO MAS32
	CLASS CORE ;
	SIZE 0.14 BY 0.16 ;
	ORIGIN 0 0 ;
	SYMMETRY X ;
	SITE core 0 0 N DO 1 BY 1 STEP 0 0 ;
	PIN P1
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0693 0.0792 0.0707 0.0808 ;
		END
	END P1
	PIN P2
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0693 0.0792 0.0707 0.0808 ;
		END
	END P2
	PIN P3
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0693 0.0792 0.0707 0.0808 ;
		END
	END P3
	PIN P4
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0693 0.0792 0.0707 0.0808 ;
		END
	END P4
	PIN P5
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0693 0.0792 0.0707 0.0808 ;
		END
	END P5
	PIN P6
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0693 0.0792 0.0707 0.0808 ;
		END
	END P6
	PIN P7
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0693 0.0792 0.0707 0.0808 ;
		END
	END P7
END MAS32

MACRO MAS33
	CLASS CORE ;
	SIZE 0.14 BY 0.16 ;
	ORIGIN 0 0 ;
	SYMMETRY X ;
	SITE core 0 0 N DO 1 BY 1 STEP 0 0 ;
	PIN P1
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0693 0.0792 0.0707 0.0808 ;
		END
	END P1
	PIN P2
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0693 0.0792 0.0707 0.0808 ;
		END
	END P2
	PIN P3
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0693 0.0792 0.0707 0.0808 ;
		END
	END P3
	PIN P4
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0693 0.0792 0.0707 0.0808 ;
		END
	END P4
	PIN P5
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0693 0.0792 0.0707 0.0808 ;
		END
	END P5
	PIN P6
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0693 0.0792 0.0707 0.0808 ;
		END
	END P6
	PIN P7
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0693 0.0792 0.0707 0.0808 ;
		END
	END P7
	PIN P8
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0693 0.0792 0.0707 0.0808 ;
		END
	END P8
END MAS33

MACRO MAS34
	CLASS CORE ;
	SIZE 0.14 BY 0.16 ;
	ORIGIN 0 0 ;
	SYMMETRY X ;
	SITE core 0 0 N DO 1 BY 1 STEP 0 0 ;
	PIN P1
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0693 0.0792 0.0707 0.0808 ;
		END
	END P1
	PIN P2
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0693 0.0792 0.0707 0.0808 ;
		END
	END P2
	PIN P3
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0693 0.0792 0.0707 0.0808 ;
		END
	END P3
	PIN P4
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0693 0.0792 0.0707 0.0808 ;
		END
	END P4
	PIN P5
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0693 0.0792 0.0707 0.0808 ;
		END
	END P5
	PIN P6
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0693 0.0792 0.0707 0.0808 ;
		END
	END P6
	PIN P7
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0693 0.0792 0.0707 0.0808 ;
		END
	END P7
	PIN P8
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0693 0.0792 0.0707 0.0808 ;
		END
	END P8
	PIN P9
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0693 0.0792 0.0707 0.0808 ;
		END
	END P9
END MAS34

MACRO MAS35
	CLASS CORE ;
	SIZE 0.16 BY 0.16 ;
	ORIGIN 0 0 ;
	SYMMETRY X ;
	SITE core 0 0 N DO 1 BY 1 STEP 0 0 ;
	PIN P1
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0792 0.0792 0.0808 0.0808 ;
		END
	END P1
	PIN P2
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0792 0.0792 0.0808 0.0808 ;
		END
	END P2
END MAS35

MACRO MAS36
	CLASS CORE ;
	SIZE 0.16 BY 0.16 ;
	ORIGIN 0 0 ;
	SYMMETRY X ;
	SITE core 0 0 N DO 1 BY 1 STEP 0 0 ;
	PIN P1
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0792 0.0792 0.0808 0.0808 ;
		END
	END P1
	PIN P2
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0792 0.0792 0.0808 0.0808 ;
		END
	END P2
	PIN P3
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0792 0.0792 0.0808 0.0808 ;
		END
	END P3
	PIN P4
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0792 0.0792 0.0808 0.0808 ;
		END
	END P4
END MAS36

MACRO MAS37
	CLASS CORE ;
	SIZE 0.16 BY 0.16 ;
	ORIGIN 0 0 ;
	SYMMETRY X ;
	SITE core 0 0 N DO 1 BY 1 STEP 0 0 ;
	PIN P1
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0792 0.0792 0.0808 0.0808 ;
		END
	END P1
	PIN P2
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0792 0.0792 0.0808 0.0808 ;
		END
	END P2
	PIN P3
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0792 0.0792 0.0808 0.0808 ;
		END
	END P3
	PIN P4
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0792 0.0792 0.0808 0.0808 ;
		END
	END P4
	PIN P5
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0792 0.0792 0.0808 0.0808 ;
		END
	END P5
END MAS37

MACRO MAS38
	CLASS CORE ;
	SIZE 0.16 BY 0.16 ;
	ORIGIN 0 0 ;
	SYMMETRY X ;
	SITE core 0 0 N DO 1 BY 1 STEP 0 0 ;
	PIN P1
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0792 0.0792 0.0808 0.0808 ;
		END
	END P1
	PIN P2
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0792 0.0792 0.0808 0.0808 ;
		END
	END P2
	PIN P3
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0792 0.0792 0.0808 0.0808 ;
		END
	END P3
	PIN P4
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0792 0.0792 0.0808 0.0808 ;
		END
	END P4
	PIN P5
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0792 0.0792 0.0808 0.0808 ;
		END
	END P5
	PIN P6
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0792 0.0792 0.0808 0.0808 ;
		END
	END P6
END MAS38

MACRO MAS39
	CLASS CORE ;
	SIZE 0.16 BY 0.16 ;
	ORIGIN 0 0 ;
	SYMMETRY X ;
	SITE core 0 0 N DO 1 BY 1 STEP 0 0 ;
	PIN P1
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0792 0.0792 0.0808 0.0808 ;
		END
	END P1
	PIN P2
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0792 0.0792 0.0808 0.0808 ;
		END
	END P2
	PIN P3
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0792 0.0792 0.0808 0.0808 ;
		END
	END P3
	PIN P4
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0792 0.0792 0.0808 0.0808 ;
		END
	END P4
	PIN P5
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0792 0.0792 0.0808 0.0808 ;
		END
	END P5
	PIN P6
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0792 0.0792 0.0808 0.0808 ;
		END
	END P6
	PIN P7
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0792 0.0792 0.0808 0.0808 ;
		END
	END P7
END MAS39

MACRO MAS40
	CLASS CORE ;
	SIZE 0.16 BY 0.16 ;
	ORIGIN 0 0 ;
	SYMMETRY X ;
	SITE core 0 0 N DO 1 BY 1 STEP 0 0 ;
	PIN P1
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0792 0.0792 0.0808 0.0808 ;
		END
	END P1
	PIN P2
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0792 0.0792 0.0808 0.0808 ;
		END
	END P2
	PIN P3
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0792 0.0792 0.0808 0.0808 ;
		END
	END P3
	PIN P4
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0792 0.0792 0.0808 0.0808 ;
		END
	END P4
	PIN P5
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0792 0.0792 0.0808 0.0808 ;
		END
	END P5
	PIN P6
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0792 0.0792 0.0808 0.0808 ;
		END
	END P6
	PIN P7
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0792 0.0792 0.0808 0.0808 ;
		END
	END P7
	PIN P8
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0792 0.0792 0.0808 0.0808 ;
		END
	END P8
END MAS40

MACRO MAS41
	CLASS CORE ;
	SIZE 0.16 BY 0.16 ;
	ORIGIN 0 0 ;
	SYMMETRY X ;
	SITE core 0 0 N DO 1 BY 1 STEP 0 0 ;
	PIN P1
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0792 0.0792 0.0808 0.0808 ;
		END
	END P1
	PIN P2
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0792 0.0792 0.0808 0.0808 ;
		END
	END P2
	PIN P3
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0792 0.0792 0.0808 0.0808 ;
		END
	END P3
	PIN P4
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0792 0.0792 0.0808 0.0808 ;
		END
	END P4
	PIN P5
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0792 0.0792 0.0808 0.0808 ;
		END
	END P5
	PIN P6
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0792 0.0792 0.0808 0.0808 ;
		END
	END P6
	PIN P7
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0792 0.0792 0.0808 0.0808 ;
		END
	END P7
	PIN P8
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0792 0.0792 0.0808 0.0808 ;
		END
	END P8
	PIN P9
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0792 0.0792 0.0808 0.0808 ;
		END
	END P9
END MAS41

MACRO MAS42
	CLASS CORE ;
	SIZE 0.18 BY 0.16 ;
	ORIGIN 0 0 ;
	SYMMETRY X ;
	SITE core 0 0 N DO 1 BY 1 STEP 0 0 ;
	PIN P1
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0891 0.0792 0.0909 0.0808 ;
		END
	END P1
	PIN P2
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0891 0.0792 0.0909 0.0808 ;
		END
	END P2
	PIN P3
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0891 0.0792 0.0909 0.0808 ;
		END
	END P3
	PIN P4
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0891 0.0792 0.0909 0.0808 ;
		END
	END P4
	PIN P5
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0891 0.0792 0.0909 0.0808 ;
		END
	END P5
END MAS42

MACRO MAS43
	CLASS CORE ;
	SIZE 0.18 BY 0.16 ;
	ORIGIN 0 0 ;
	SYMMETRY X ;
	SITE core 0 0 N DO 1 BY 1 STEP 0 0 ;
	PIN P1
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0891 0.0792 0.0909 0.0808 ;
		END
	END P1
	PIN P2
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0891 0.0792 0.0909 0.0808 ;
		END
	END P2
	PIN P3
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0891 0.0792 0.0909 0.0808 ;
		END
	END P3
	PIN P4
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0891 0.0792 0.0909 0.0808 ;
		END
	END P4
	PIN P5
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0891 0.0792 0.0909 0.0808 ;
		END
	END P5
	PIN P6
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0891 0.0792 0.0909 0.0808 ;
		END
	END P6
END MAS43

MACRO MAS44
	CLASS CORE ;
	SIZE 0.18 BY 0.16 ;
	ORIGIN 0 0 ;
	SYMMETRY X ;
	SITE core 0 0 N DO 1 BY 1 STEP 0 0 ;
	PIN P1
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0891 0.0792 0.0909 0.0808 ;
		END
	END P1
	PIN P2
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0891 0.0792 0.0909 0.0808 ;
		END
	END P2
	PIN P3
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0891 0.0792 0.0909 0.0808 ;
		END
	END P3
	PIN P4
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0891 0.0792 0.0909 0.0808 ;
		END
	END P4
	PIN P5
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0891 0.0792 0.0909 0.0808 ;
		END
	END P5
	PIN P6
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0891 0.0792 0.0909 0.0808 ;
		END
	END P6
	PIN P7
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0891 0.0792 0.0909 0.0808 ;
		END
	END P7
END MAS44

MACRO MAS45
	CLASS CORE ;
	SIZE 0.18 BY 0.16 ;
	ORIGIN 0 0 ;
	SYMMETRY X ;
	SITE core 0 0 N DO 1 BY 1 STEP 0 0 ;
	PIN P1
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0891 0.0792 0.0909 0.0808 ;
		END
	END P1
	PIN P2
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0891 0.0792 0.0909 0.0808 ;
		END
	END P2
	PIN P3
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0891 0.0792 0.0909 0.0808 ;
		END
	END P3
	PIN P4
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0891 0.0792 0.0909 0.0808 ;
		END
	END P4
	PIN P5
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0891 0.0792 0.0909 0.0808 ;
		END
	END P5
	PIN P6
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0891 0.0792 0.0909 0.0808 ;
		END
	END P6
	PIN P7
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0891 0.0792 0.0909 0.0808 ;
		END
	END P7
	PIN P8
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0891 0.0792 0.0909 0.0808 ;
		END
	END P8
	PIN P9
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.0891 0.0792 0.0909 0.0808 ;
		END
	END P9
END MAS45

MACRO MAS46
	CLASS CORE ;
	SIZE 0.2 BY 0.16 ;
	ORIGIN 0 0 ;
	SYMMETRY X ;
	SITE core 0 0 N DO 1 BY 1 STEP 0 0 ;
	PIN P1
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.099 0.0792 0.101 0.0808 ;
		END
	END P1
	PIN P2
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.099 0.0792 0.101 0.0808 ;
		END
	END P2
END MAS46

MACRO MAS47
	CLASS CORE ;
	SIZE 0.2 BY 0.16 ;
	ORIGIN 0 0 ;
	SYMMETRY X ;
	SITE core 0 0 N DO 1 BY 1 STEP 0 0 ;
	PIN P1
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.099 0.0792 0.101 0.0808 ;
		END
	END P1
	PIN P2
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.099 0.0792 0.101 0.0808 ;
		END
	END P2
	PIN P3
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.099 0.0792 0.101 0.0808 ;
		END
	END P3
	PIN P4
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.099 0.0792 0.101 0.0808 ;
		END
	END P4
END MAS47

MACRO MAS48
	CLASS CORE ;
	SIZE 0.2 BY 0.16 ;
	ORIGIN 0 0 ;
	SYMMETRY X ;
	SITE core 0 0 N DO 1 BY 1 STEP 0 0 ;
	PIN P1
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.099 0.0792 0.101 0.0808 ;
		END
	END P1
	PIN P2
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.099 0.0792 0.101 0.0808 ;
		END
	END P2
	PIN P3
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.099 0.0792 0.101 0.0808 ;
		END
	END P3
	PIN P4
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.099 0.0792 0.101 0.0808 ;
		END
	END P4
	PIN P5
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.099 0.0792 0.101 0.0808 ;
		END
	END P5
END MAS48

MACRO MAS49
	CLASS CORE ;
	SIZE 0.2 BY 0.16 ;
	ORIGIN 0 0 ;
	SYMMETRY X ;
	SITE core 0 0 N DO 1 BY 1 STEP 0 0 ;
	PIN P1
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.099 0.0792 0.101 0.0808 ;
		END
	END P1
	PIN P2
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.099 0.0792 0.101 0.0808 ;
		END
	END P2
	PIN P3
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.099 0.0792 0.101 0.0808 ;
		END
	END P3
	PIN P4
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.099 0.0792 0.101 0.0808 ;
		END
	END P4
	PIN P5
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.099 0.0792 0.101 0.0808 ;
		END
	END P5
	PIN P6
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.099 0.0792 0.101 0.0808 ;
		END
	END P6
END MAS49

MACRO MAS50
	CLASS CORE ;
	SIZE 0.24 BY 0.16 ;
	ORIGIN 0 0 ;
	SYMMETRY X ;
	SITE core 0 0 N DO 1 BY 1 STEP 0 0 ;
	PIN P1
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.1188 0.0792 0.1212 0.0808 ;
		END
	END P1
	PIN P2
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.1188 0.0792 0.1212 0.0808 ;
		END
	END P2
END MAS50

MACRO MAS51
	CLASS CORE ;
	SIZE 0.26 BY 0.16 ;
	ORIGIN 0 0 ;
	SYMMETRY X ;
	SITE core 0 0 N DO 1 BY 1 STEP 0 0 ;
	PIN P1
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.1287 0.0792 0.1313 0.0808 ;
		END
	END P1
	PIN P2
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.1287 0.0792 0.1313 0.0808 ;
		END
	END P2
	PIN P3
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.1287 0.0792 0.1313 0.0808 ;
		END
	END P3
	PIN P4
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.1287 0.0792 0.1313 0.0808 ;
		END
	END P4
	PIN P5
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.1287 0.0792 0.1313 0.0808 ;
		END
	END P5
	PIN P6
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.1287 0.0792 0.1313 0.0808 ;
		END
	END P6
	PIN P7
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.1287 0.0792 0.1313 0.0808 ;
		END
	END P7
	PIN P8
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.1287 0.0792 0.1313 0.0808 ;
		END
	END P8
	PIN P9
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.1287 0.0792 0.1313 0.0808 ;
		END
	END P9
END MAS51

MACRO MAS52
	CLASS CORE ;
	SIZE 0.28 BY 0.16 ;
	ORIGIN 0 0 ;
	SYMMETRY X ;
	SITE core 0 0 N DO 1 BY 1 STEP 0 0 ;
	PIN P1
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.1386 0.0792 0.1414 0.0808 ;
		END
	END P1
	PIN P2
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.1386 0.0792 0.1414 0.0808 ;
		END
	END P2
	PIN P3
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.1386 0.0792 0.1414 0.0808 ;
		END
	END P3
	PIN P4
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.1386 0.0792 0.1414 0.0808 ;
		END
	END P4
	PIN P5
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.1386 0.0792 0.1414 0.0808 ;
		END
	END P5
	PIN P6
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.1386 0.0792 0.1414 0.0808 ;
		END
	END P6
	PIN P7
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.1386 0.0792 0.1414 0.0808 ;
		END
	END P7
	PIN P8
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.1386 0.0792 0.1414 0.0808 ;
		END
	END P8
	PIN P9
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.1386 0.0792 0.1414 0.0808 ;
		END
	END P9
END MAS52

MACRO MAS53
	CLASS CORE ;
	SIZE 0.32 BY 0.16 ;
	ORIGIN 0 0 ;
	SYMMETRY X ;
	SITE core 0 0 N DO 1 BY 1 STEP 0 0 ;
	PIN P1
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.1584 0.0792 0.1616 0.0808 ;
		END
	END P1
	PIN P2
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.1584 0.0792 0.1616 0.0808 ;
		END
	END P2
	PIN P3
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.1584 0.0792 0.1616 0.0808 ;
		END
	END P3
END MAS53

MACRO MAS54
	CLASS CORE ;
	SIZE 0.4 BY 0.16 ;
	ORIGIN 0 0 ;
	SYMMETRY X ;
	SITE core 0 0 N DO 1 BY 1 STEP 0 0 ;
	PIN P1
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.198 0.0792 0.202 0.0808 ;
		END
	END P1
	PIN P2
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.198 0.0792 0.202 0.0808 ;
		END
	END P2
	PIN P3
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.198 0.0792 0.202 0.0808 ;
		END
	END P3
END MAS54

MACRO MAS55
	CLASS CORE ;
	SIZE 1 BY 0.16 ;
	ORIGIN 0 0 ;
	SYMMETRY X ;
	SITE core 0 0 N DO 1 BY 1 STEP 0 0 ;
	PIN P1
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.495 0.0792 0.505 0.0808 ;
		END
	END P1
	PIN P2
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.495 0.0792 0.505 0.0808 ;
		END
	END P2
END MAS55

MACRO MAS56
	CLASS CORE ;
	SIZE 0.8 BY 0.96 ;
	ORIGIN 0 0 ;
	SYMMETRY X ;
	SITE core 0 0 N DO 1 BY 1 STEP 0 0 ;
	PIN P1
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.396 0.4752 0.404 0.4848 ;
		END
	END P1
	PIN P2
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.396 0.4752 0.404 0.4848 ;
		END
	END P2
END MAS56

MACRO MAS57
	CLASS CORE ;
	SIZE 0.8 BY 0.96 ;
	ORIGIN 0 0 ;
	SYMMETRY X ;
	SITE core 0 0 N DO 1 BY 1 STEP 0 0 ;
	PIN P1
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.396 0.4752 0.404 0.4848 ;
		END
	END P1
	PIN P2
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.396 0.4752 0.404 0.4848 ;
		END
	END P2
	PIN P3
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.396 0.4752 0.404 0.4848 ;
		END
	END P3
END MAS57

MACRO MAS58
	CLASS CORE ;
	SIZE 0.8 BY 0.96 ;
	ORIGIN 0 0 ;
	SYMMETRY X ;
	SITE core 0 0 N DO 1 BY 1 STEP 0 0 ;
	PIN P1
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.396 0.4752 0.404 0.4848 ;
		END
	END P1
	PIN P2
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.396 0.4752 0.404 0.4848 ;
		END
	END P2
	PIN P3
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.396 0.4752 0.404 0.4848 ;
		END
	END P3
	PIN P4
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.396 0.4752 0.404 0.4848 ;
		END
	END P4
END MAS58

MACRO MAS59
	CLASS CORE ;
	SIZE 0.8 BY 0.96 ;
	ORIGIN 0 0 ;
	SYMMETRY X ;
	SITE core 0 0 N DO 1 BY 1 STEP 0 0 ;
	PIN P1
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.396 0.4752 0.404 0.4848 ;
		END
	END P1
	PIN P2
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.396 0.4752 0.404 0.4848 ;
		END
	END P2
	PIN P3
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.396 0.4752 0.404 0.4848 ;
		END
	END P3
	PIN P4
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.396 0.4752 0.404 0.4848 ;
		END
	END P4
	PIN P5
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.396 0.4752 0.404 0.4848 ;
		END
	END P5
END MAS59

MACRO MAS60
	CLASS CORE ;
	SIZE 0.8 BY 0.96 ;
	ORIGIN 0 0 ;
	SYMMETRY X ;
	SITE core 0 0 N DO 1 BY 1 STEP 0 0 ;
	PIN P1
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.396 0.4752 0.404 0.4848 ;
		END
	END P1
	PIN P2
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.396 0.4752 0.404 0.4848 ;
		END
	END P2
	PIN P3
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.396 0.4752 0.404 0.4848 ;
		END
	END P3
	PIN P4
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.396 0.4752 0.404 0.4848 ;
		END
	END P4
	PIN P5
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.396 0.4752 0.404 0.4848 ;
		END
	END P5
	PIN P6
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.396 0.4752 0.404 0.4848 ;
		END
	END P6
END MAS60

MACRO MAS61
	CLASS CORE ;
	SIZE 0.8 BY 0.96 ;
	ORIGIN 0 0 ;
	SYMMETRY X ;
	SITE core 0 0 N DO 1 BY 1 STEP 0 0 ;
	PIN P1
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.396 0.4752 0.404 0.4848 ;
		END
	END P1
	PIN P2
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.396 0.4752 0.404 0.4848 ;
		END
	END P2
	PIN P3
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.396 0.4752 0.404 0.4848 ;
		END
	END P3
	PIN P4
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.396 0.4752 0.404 0.4848 ;
		END
	END P4
	PIN P5
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.396 0.4752 0.404 0.4848 ;
		END
	END P5
	PIN P6
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.396 0.4752 0.404 0.4848 ;
		END
	END P6
	PIN P7
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.396 0.4752 0.404 0.4848 ;
		END
	END P7
END MAS61

MACRO MAS62
	CLASS CORE ;
	SIZE 0.8 BY 0.96 ;
	ORIGIN 0 0 ;
	SYMMETRY X ;
	SITE core 0 0 N DO 1 BY 1 STEP 0 0 ;
	PIN P1
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.396 0.4752 0.404 0.4848 ;
		END
	END P1
	PIN P2
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.396 0.4752 0.404 0.4848 ;
		END
	END P2
	PIN P3
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.396 0.4752 0.404 0.4848 ;
		END
	END P3
	PIN P4
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.396 0.4752 0.404 0.4848 ;
		END
	END P4
	PIN P5
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.396 0.4752 0.404 0.4848 ;
		END
	END P5
	PIN P6
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.396 0.4752 0.404 0.4848 ;
		END
	END P6
	PIN P7
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.396 0.4752 0.404 0.4848 ;
		END
	END P7
	PIN P8
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 0.396 0.4752 0.404 0.4848 ;
		END
	END P8
END MAS62

MACRO MAS63
	CLASS CORE ;
	SIZE 2.79 BY 2.88 ;
	ORIGIN 0 0 ;
	SYMMETRY X ;
	SITE core 0 0 N DO 1 BY 1 STEP 0 0 ;
	PIN P1
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 1.38105 1.4256 1.40895 1.4544 ;
		END
	END P1
	PIN P2
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 1.38105 1.4256 1.40895 1.4544 ;
		END
	END P2
	PIN P3
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 1.38105 1.4256 1.40895 1.4544 ;
		END
	END P3
	PIN P4
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 1.38105 1.4256 1.40895 1.4544 ;
		END
	END P4
	PIN P5
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 1.38105 1.4256 1.40895 1.4544 ;
		END
	END P5
	PIN P6
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 1.38105 1.4256 1.40895 1.4544 ;
		END
	END P6
	PIN P7
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 1.38105 1.4256 1.40895 1.4544 ;
		END
	END P7
	PIN P8
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 1.38105 1.4256 1.40895 1.4544 ;
		END
	END P8
	PIN P9
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 1.38105 1.4256 1.40895 1.4544 ;
		END
	END P9
	PIN P10
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 1.38105 1.4256 1.40895 1.4544 ;
		END
	END P10
	PIN P11
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 1.38105 1.4256 1.40895 1.4544 ;
		END
	END P11
	PIN P12
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 1.38105 1.4256 1.40895 1.4544 ;
		END
	END P12
	PIN P13
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 1.38105 1.4256 1.40895 1.4544 ;
		END
	END P13
	PIN P14
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 1.38105 1.4256 1.40895 1.4544 ;
		END
	END P14
	PIN P15
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 1.38105 1.4256 1.40895 1.4544 ;
		END
	END P15
	PIN P16
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 1.38105 1.4256 1.40895 1.4544 ;
		END
	END P16
	PIN P17
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 1.38105 1.4256 1.40895 1.4544 ;
		END
	END P17
	PIN P18
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 1.38105 1.4256 1.40895 1.4544 ;
		END
	END P18
	PIN P19
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 1.38105 1.4256 1.40895 1.4544 ;
		END
	END P19
	PIN P20
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 1.38105 1.4256 1.40895 1.4544 ;
		END
	END P20
	PIN P21
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 1.38105 1.4256 1.40895 1.4544 ;
		END
	END P21
	PIN P22
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 1.38105 1.4256 1.40895 1.4544 ;
		END
	END P22
	PIN P23
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 1.38105 1.4256 1.40895 1.4544 ;
		END
	END P23
	PIN P24
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 1.38105 1.4256 1.40895 1.4544 ;
		END
	END P24
	PIN P25
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 1.38105 1.4256 1.40895 1.4544 ;
		END
	END P25
	PIN P26
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 1.38105 1.4256 1.40895 1.4544 ;
		END
	END P26
	PIN P27
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 1.38105 1.4256 1.40895 1.4544 ;
		END
	END P27
	PIN P28
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 1.38105 1.4256 1.40895 1.4544 ;
		END
	END P28
	PIN P29
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 1.38105 1.4256 1.40895 1.4544 ;
		END
	END P29
END MAS63

MACRO MAS64
	CLASS CORE ;
	SIZE 2.79 BY 2.88 ;
	ORIGIN 0 0 ;
	SYMMETRY X ;
	SITE core 0 0 N DO 1 BY 1 STEP 0 0 ;
	PIN P1
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 1.38105 1.4256 1.40895 1.4544 ;
		END
	END P1
	PIN P2
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 1.38105 1.4256 1.40895 1.4544 ;
		END
	END P2
	PIN P3
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 1.38105 1.4256 1.40895 1.4544 ;
		END
	END P3
	PIN P4
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 1.38105 1.4256 1.40895 1.4544 ;
		END
	END P4
	PIN P5
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 1.38105 1.4256 1.40895 1.4544 ;
		END
	END P5
	PIN P6
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 1.38105 1.4256 1.40895 1.4544 ;
		END
	END P6
	PIN P7
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 1.38105 1.4256 1.40895 1.4544 ;
		END
	END P7
	PIN P8
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 1.38105 1.4256 1.40895 1.4544 ;
		END
	END P8
	PIN P9
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 1.38105 1.4256 1.40895 1.4544 ;
		END
	END P9
	PIN P10
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 1.38105 1.4256 1.40895 1.4544 ;
		END
	END P10
	PIN P11
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 1.38105 1.4256 1.40895 1.4544 ;
		END
	END P11
	PIN P12
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 1.38105 1.4256 1.40895 1.4544 ;
		END
	END P12
	PIN P13
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 1.38105 1.4256 1.40895 1.4544 ;
		END
	END P13
	PIN P14
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 1.38105 1.4256 1.40895 1.4544 ;
		END
	END P14
	PIN P15
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 1.38105 1.4256 1.40895 1.4544 ;
		END
	END P15
	PIN P16
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 1.38105 1.4256 1.40895 1.4544 ;
		END
	END P16
	PIN P17
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 1.38105 1.4256 1.40895 1.4544 ;
		END
	END P17
	PIN P18
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 1.38105 1.4256 1.40895 1.4544 ;
		END
	END P18
	PIN P19
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 1.38105 1.4256 1.40895 1.4544 ;
		END
	END P19
	PIN P20
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 1.38105 1.4256 1.40895 1.4544 ;
		END
	END P20
	PIN P21
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 1.38105 1.4256 1.40895 1.4544 ;
		END
	END P21
	PIN P22
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 1.38105 1.4256 1.40895 1.4544 ;
		END
	END P22
	PIN P23
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 1.38105 1.4256 1.40895 1.4544 ;
		END
	END P23
	PIN P24
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 1.38105 1.4256 1.40895 1.4544 ;
		END
	END P24
	PIN P25
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 1.38105 1.4256 1.40895 1.4544 ;
		END
	END P25
	PIN P26
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 1.38105 1.4256 1.40895 1.4544 ;
		END
	END P26
	PIN P27
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 1.38105 1.4256 1.40895 1.4544 ;
		END
	END P27
	PIN P28
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 1.38105 1.4256 1.40895 1.4544 ;
		END
	END P28
	PIN P29
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 1.38105 1.4256 1.40895 1.4544 ;
		END
	END P29
	PIN P30
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 1.38105 1.4256 1.40895 1.4544 ;
		END
	END P30
	PIN P31
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 1.38105 1.4256 1.40895 1.4544 ;
		END
	END P31
	PIN P32
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 1.38105 1.4256 1.40895 1.4544 ;
		END
	END P32
END MAS64

MACRO MAS65
	CLASS CORE ;
	SIZE 3.68 BY 3.68 ;
	ORIGIN 0 0 ;
	SYMMETRY X ;
	SITE core 0 0 N DO 1 BY 1 STEP 0 0 ;
	PIN P1
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 1.8216 1.8216 1.8584 1.8584 ;
		END
	END P1
	PIN P2
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 1.8216 1.8216 1.8584 1.8584 ;
		END
	END P2
	PIN P3
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 1.8216 1.8216 1.8584 1.8584 ;
		END
	END P3
	PIN P4
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 1.8216 1.8216 1.8584 1.8584 ;
		END
	END P4
	PIN P5
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 1.8216 1.8216 1.8584 1.8584 ;
		END
	END P5
	PIN P6
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 1.8216 1.8216 1.8584 1.8584 ;
		END
	END P6
	PIN P7
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 1.8216 1.8216 1.8584 1.8584 ;
		END
	END P7
	PIN P8
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 1.8216 1.8216 1.8584 1.8584 ;
		END
	END P8
	PIN P9
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 1.8216 1.8216 1.8584 1.8584 ;
		END
	END P9
	PIN P10
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 1.8216 1.8216 1.8584 1.8584 ;
		END
	END P10
	PIN P11
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 1.8216 1.8216 1.8584 1.8584 ;
		END
	END P11
	PIN P12
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 1.8216 1.8216 1.8584 1.8584 ;
		END
	END P12
	PIN P13
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 1.8216 1.8216 1.8584 1.8584 ;
		END
	END P13
	PIN P14
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 1.8216 1.8216 1.8584 1.8584 ;
		END
	END P14
	PIN P15
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 1.8216 1.8216 1.8584 1.8584 ;
		END
	END P15
	PIN P16
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 1.8216 1.8216 1.8584 1.8584 ;
		END
	END P16
	PIN P17
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 1.8216 1.8216 1.8584 1.8584 ;
		END
	END P17
	PIN P18
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 1.8216 1.8216 1.8584 1.8584 ;
		END
	END P18
	PIN P19
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 1.8216 1.8216 1.8584 1.8584 ;
		END
	END P19
	PIN P20
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 1.8216 1.8216 1.8584 1.8584 ;
		END
	END P20
	PIN P21
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 1.8216 1.8216 1.8584 1.8584 ;
		END
	END P21
	PIN P22
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 1.8216 1.8216 1.8584 1.8584 ;
		END
	END P22
	PIN P23
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 1.8216 1.8216 1.8584 1.8584 ;
		END
	END P23
	PIN P24
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 1.8216 1.8216 1.8584 1.8584 ;
		END
	END P24
	PIN P25
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 1.8216 1.8216 1.8584 1.8584 ;
		END
	END P25
	PIN P26
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 1.8216 1.8216 1.8584 1.8584 ;
		END
	END P26
	PIN P27
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 1.8216 1.8216 1.8584 1.8584 ;
		END
	END P27
	PIN P28
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 1.8216 1.8216 1.8584 1.8584 ;
		END
	END P28
	PIN P29
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 1.8216 1.8216 1.8584 1.8584 ;
		END
	END P29
	PIN P30
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 1.8216 1.8216 1.8584 1.8584 ;
		END
	END P30
	PIN P31
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 1.8216 1.8216 1.8584 1.8584 ;
		END
	END P31
	PIN P32
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 1.8216 1.8216 1.8584 1.8584 ;
		END
	END P32
	PIN P33
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 1.8216 1.8216 1.8584 1.8584 ;
		END
	END P33
	PIN P34
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 1.8216 1.8216 1.8584 1.8584 ;
		END
	END P34
	PIN P35
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 1.8216 1.8216 1.8584 1.8584 ;
		END
	END P35
	PIN P36
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 1.8216 1.8216 1.8584 1.8584 ;
		END
	END P36
	PIN P37
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 1.8216 1.8216 1.8584 1.8584 ;
		END
	END P37
	PIN P38
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 1.8216 1.8216 1.8584 1.8584 ;
		END
	END P38
	PIN P39
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 1.8216 1.8216 1.8584 1.8584 ;
		END
	END P39
	PIN P40
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 1.8216 1.8216 1.8584 1.8584 ;
		END
	END P40
	PIN P41
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 1.8216 1.8216 1.8584 1.8584 ;
		END
	END P41
	PIN P42
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 1.8216 1.8216 1.8584 1.8584 ;
		END
	END P42
	PIN P43
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 1.8216 1.8216 1.8584 1.8584 ;
		END
	END P43
	PIN P44
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 1.8216 1.8216 1.8584 1.8584 ;
		END
	END P44
	PIN P45
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 1.8216 1.8216 1.8584 1.8584 ;
		END
	END P45
	PIN P46
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 1.8216 1.8216 1.8584 1.8584 ;
		END
	END P46
	PIN P47
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 1.8216 1.8216 1.8584 1.8584 ;
		END
	END P47
	PIN P48
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 1.8216 1.8216 1.8584 1.8584 ;
		END
	END P48
	PIN P49
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 1.8216 1.8216 1.8584 1.8584 ;
		END
	END P49
	PIN P50
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 1.8216 1.8216 1.8584 1.8584 ;
		END
	END P50
	PIN P51
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 1.8216 1.8216 1.8584 1.8584 ;
		END
	END P51
END MAS65

MACRO MAS66
	CLASS CORE ;
	SIZE 5.24 BY 5.28 ;
	ORIGIN 0 0 ;
	SYMMETRY X ;
	SITE core 0 0 N DO 1 BY 1 STEP 0 0 ;
	PIN P1
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 2.5938 2.6136 2.6462 2.6664 ;
		END
	END P1
	PIN P2
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 2.5938 2.6136 2.6462 2.6664 ;
		END
	END P2
	PIN P3
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 2.5938 2.6136 2.6462 2.6664 ;
		END
	END P3
	PIN P4
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 2.5938 2.6136 2.6462 2.6664 ;
		END
	END P4
	PIN P5
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 2.5938 2.6136 2.6462 2.6664 ;
		END
	END P5
	PIN P6
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 2.5938 2.6136 2.6462 2.6664 ;
		END
	END P6
	PIN P7
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 2.5938 2.6136 2.6462 2.6664 ;
		END
	END P7
	PIN P8
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 2.5938 2.6136 2.6462 2.6664 ;
		END
	END P8
	PIN P9
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 2.5938 2.6136 2.6462 2.6664 ;
		END
	END P9
	PIN P10
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 2.5938 2.6136 2.6462 2.6664 ;
		END
	END P10
	PIN P11
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 2.5938 2.6136 2.6462 2.6664 ;
		END
	END P11
	PIN P12
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 2.5938 2.6136 2.6462 2.6664 ;
		END
	END P12
	PIN P13
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 2.5938 2.6136 2.6462 2.6664 ;
		END
	END P13
	PIN P14
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 2.5938 2.6136 2.6462 2.6664 ;
		END
	END P14
	PIN P15
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 2.5938 2.6136 2.6462 2.6664 ;
		END
	END P15
	PIN P16
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 2.5938 2.6136 2.6462 2.6664 ;
		END
	END P16
	PIN P17
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 2.5938 2.6136 2.6462 2.6664 ;
		END
	END P17
	PIN P18
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 2.5938 2.6136 2.6462 2.6664 ;
		END
	END P18
	PIN P19
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 2.5938 2.6136 2.6462 2.6664 ;
		END
	END P19
	PIN P20
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 2.5938 2.6136 2.6462 2.6664 ;
		END
	END P20
	PIN P21
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 2.5938 2.6136 2.6462 2.6664 ;
		END
	END P21
	PIN P22
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 2.5938 2.6136 2.6462 2.6664 ;
		END
	END P22
	PIN P23
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 2.5938 2.6136 2.6462 2.6664 ;
		END
	END P23
	PIN P24
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 2.5938 2.6136 2.6462 2.6664 ;
		END
	END P24
	PIN P25
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 2.5938 2.6136 2.6462 2.6664 ;
		END
	END P25
	PIN P26
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 2.5938 2.6136 2.6462 2.6664 ;
		END
	END P26
	PIN P27
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 2.5938 2.6136 2.6462 2.6664 ;
		END
	END P27
	PIN P28
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 2.5938 2.6136 2.6462 2.6664 ;
		END
	END P28
	PIN P29
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 2.5938 2.6136 2.6462 2.6664 ;
		END
	END P29
	PIN P30
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 2.5938 2.6136 2.6462 2.6664 ;
		END
	END P30
	PIN P31
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 2.5938 2.6136 2.6462 2.6664 ;
		END
	END P31
	PIN P32
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 2.5938 2.6136 2.6462 2.6664 ;
		END
	END P32
	PIN P33
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 2.5938 2.6136 2.6462 2.6664 ;
		END
	END P33
	PIN P34
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 2.5938 2.6136 2.6462 2.6664 ;
		END
	END P34
	PIN P35
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 2.5938 2.6136 2.6462 2.6664 ;
		END
	END P35
	PIN P36
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 2.5938 2.6136 2.6462 2.6664 ;
		END
	END P36
	PIN P37
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 2.5938 2.6136 2.6462 2.6664 ;
		END
	END P37
	PIN P38
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 2.5938 2.6136 2.6462 2.6664 ;
		END
	END P38
	PIN P39
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 2.5938 2.6136 2.6462 2.6664 ;
		END
	END P39
	PIN P40
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 2.5938 2.6136 2.6462 2.6664 ;
		END
	END P40
	PIN P41
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 2.5938 2.6136 2.6462 2.6664 ;
		END
	END P41
	PIN P42
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 2.5938 2.6136 2.6462 2.6664 ;
		END
	END P42
	PIN P43
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 2.5938 2.6136 2.6462 2.6664 ;
		END
	END P43
	PIN P44
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 2.5938 2.6136 2.6462 2.6664 ;
		END
	END P44
	PIN P45
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 2.5938 2.6136 2.6462 2.6664 ;
		END
	END P45
	PIN P46
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 2.5938 2.6136 2.6462 2.6664 ;
		END
	END P46
	PIN P47
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 2.5938 2.6136 2.6462 2.6664 ;
		END
	END P47
	PIN P48
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 2.5938 2.6136 2.6462 2.6664 ;
		END
	END P48
	PIN P49
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 2.5938 2.6136 2.6462 2.6664 ;
		END
	END P49
	PIN P50
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 2.5938 2.6136 2.6462 2.6664 ;
		END
	END P50
	PIN P51
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 2.5938 2.6136 2.6462 2.6664 ;
		END
	END P51
END MAS66

MACRO MAS67
	CLASS CORE ;
	SIZE 6.52 BY 6.4 ;
	ORIGIN 0 0 ;
	SYMMETRY X ;
	SITE core 0 0 N DO 1 BY 1 STEP 0 0 ;
	PIN P1
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 3.2274 3.168 3.2926 3.232 ;
		END
	END P1
	PIN P2
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 3.2274 3.168 3.2926 3.232 ;
		END
	END P2
	PIN P3
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 3.2274 3.168 3.2926 3.232 ;
		END
	END P3
	PIN P4
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 3.2274 3.168 3.2926 3.232 ;
		END
	END P4
	PIN P5
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 3.2274 3.168 3.2926 3.232 ;
		END
	END P5
	PIN P6
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 3.2274 3.168 3.2926 3.232 ;
		END
	END P6
	PIN P7
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 3.2274 3.168 3.2926 3.232 ;
		END
	END P7
	PIN P8
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 3.2274 3.168 3.2926 3.232 ;
		END
	END P8
	PIN P9
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 3.2274 3.168 3.2926 3.232 ;
		END
	END P9
	PIN P10
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 3.2274 3.168 3.2926 3.232 ;
		END
	END P10
	PIN P11
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 3.2274 3.168 3.2926 3.232 ;
		END
	END P11
	PIN P12
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 3.2274 3.168 3.2926 3.232 ;
		END
	END P12
	PIN P13
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 3.2274 3.168 3.2926 3.232 ;
		END
	END P13
	PIN P14
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 3.2274 3.168 3.2926 3.232 ;
		END
	END P14
	PIN P15
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 3.2274 3.168 3.2926 3.232 ;
		END
	END P15
	PIN P16
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 3.2274 3.168 3.2926 3.232 ;
		END
	END P16
	PIN P17
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 3.2274 3.168 3.2926 3.232 ;
		END
	END P17
	PIN P18
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 3.2274 3.168 3.2926 3.232 ;
		END
	END P18
	PIN P19
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 3.2274 3.168 3.2926 3.232 ;
		END
	END P19
	PIN P20
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 3.2274 3.168 3.2926 3.232 ;
		END
	END P20
	PIN P21
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 3.2274 3.168 3.2926 3.232 ;
		END
	END P21
	PIN P22
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 3.2274 3.168 3.2926 3.232 ;
		END
	END P22
	PIN P23
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 3.2274 3.168 3.2926 3.232 ;
		END
	END P23
	PIN P24
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 3.2274 3.168 3.2926 3.232 ;
		END
	END P24
	PIN P25
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 3.2274 3.168 3.2926 3.232 ;
		END
	END P25
	PIN P26
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 3.2274 3.168 3.2926 3.232 ;
		END
	END P26
	PIN P27
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 3.2274 3.168 3.2926 3.232 ;
		END
	END P27
	PIN P28
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 3.2274 3.168 3.2926 3.232 ;
		END
	END P28
	PIN P29
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 3.2274 3.168 3.2926 3.232 ;
		END
	END P29
	PIN P30
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 3.2274 3.168 3.2926 3.232 ;
		END
	END P30
	PIN P31
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 3.2274 3.168 3.2926 3.232 ;
		END
	END P31
	PIN P32
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 3.2274 3.168 3.2926 3.232 ;
		END
	END P32
	PIN P33
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 3.2274 3.168 3.2926 3.232 ;
		END
	END P33
	PIN P34
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 3.2274 3.168 3.2926 3.232 ;
		END
	END P34
	PIN P35
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 3.2274 3.168 3.2926 3.232 ;
		END
	END P35
	PIN P36
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 3.2274 3.168 3.2926 3.232 ;
		END
	END P36
	PIN P37
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 3.2274 3.168 3.2926 3.232 ;
		END
	END P37
	PIN P38
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 3.2274 3.168 3.2926 3.232 ;
		END
	END P38
	PIN P39
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 3.2274 3.168 3.2926 3.232 ;
		END
	END P39
	PIN P40
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 3.2274 3.168 3.2926 3.232 ;
		END
	END P40
	PIN P41
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 3.2274 3.168 3.2926 3.232 ;
		END
	END P41
	PIN P42
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 3.2274 3.168 3.2926 3.232 ;
		END
	END P42
	PIN P43
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 3.2274 3.168 3.2926 3.232 ;
		END
	END P43
	PIN P44
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 3.2274 3.168 3.2926 3.232 ;
		END
	END P44
	PIN P45
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 3.2274 3.168 3.2926 3.232 ;
		END
	END P45
	PIN P46
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 3.2274 3.168 3.2926 3.232 ;
		END
	END P46
	PIN P47
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 3.2274 3.168 3.2926 3.232 ;
		END
	END P47
	PIN P48
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 3.2274 3.168 3.2926 3.232 ;
		END
	END P48
	PIN P49
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 3.2274 3.168 3.2926 3.232 ;
		END
	END P49
	PIN P50
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 3.2274 3.168 3.2926 3.232 ;
		END
	END P50
	PIN P51
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 3.2274 3.168 3.2926 3.232 ;
		END
	END P51
	PIN P52
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 3.2274 3.168 3.2926 3.232 ;
		END
	END P52
	PIN P53
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 3.2274 3.168 3.2926 3.232 ;
		END
	END P53
	PIN P54
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 3.2274 3.168 3.2926 3.232 ;
		END
	END P54
	PIN P55
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 3.2274 3.168 3.2926 3.232 ;
		END
	END P55
	PIN P56
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 3.2274 3.168 3.2926 3.232 ;
		END
	END P56
	PIN P57
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 3.2274 3.168 3.2926 3.232 ;
		END
	END P57
	PIN P58
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 3.2274 3.168 3.2926 3.232 ;
		END
	END P58
	PIN P59
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 3.2274 3.168 3.2926 3.232 ;
		END
	END P59
	PIN P60
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 3.2274 3.168 3.2926 3.232 ;
		END
	END P60
END MAS67

MACRO MAS68
	CLASS CORE ;
	SIZE 7.21 BY 7.2 ;
	ORIGIN 0 0 ;
	SYMMETRY X ;
	SITE core 0 0 N DO 1 BY 1 STEP 0 0 ;
	PIN P1
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 3.56895 3.564 3.64105 3.636 ;
		END
	END P1
	PIN P2
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 3.56895 3.564 3.64105 3.636 ;
		END
	END P2
	PIN P3
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 3.56895 3.564 3.64105 3.636 ;
		END
	END P3
	PIN P4
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 3.56895 3.564 3.64105 3.636 ;
		END
	END P4
	PIN P5
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 3.56895 3.564 3.64105 3.636 ;
		END
	END P5
	PIN P6
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 3.56895 3.564 3.64105 3.636 ;
		END
	END P6
	PIN P7
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 3.56895 3.564 3.64105 3.636 ;
		END
	END P7
	PIN P8
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 3.56895 3.564 3.64105 3.636 ;
		END
	END P8
	PIN P9
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 3.56895 3.564 3.64105 3.636 ;
		END
	END P9
	PIN P10
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 3.56895 3.564 3.64105 3.636 ;
		END
	END P10
	PIN P11
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 3.56895 3.564 3.64105 3.636 ;
		END
	END P11
	PIN P12
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 3.56895 3.564 3.64105 3.636 ;
		END
	END P12
	PIN P13
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 3.56895 3.564 3.64105 3.636 ;
		END
	END P13
	PIN P14
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 3.56895 3.564 3.64105 3.636 ;
		END
	END P14
	PIN P15
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 3.56895 3.564 3.64105 3.636 ;
		END
	END P15
	PIN P16
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 3.56895 3.564 3.64105 3.636 ;
		END
	END P16
	PIN P17
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 3.56895 3.564 3.64105 3.636 ;
		END
	END P17
	PIN P18
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 3.56895 3.564 3.64105 3.636 ;
		END
	END P18
	PIN P19
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 3.56895 3.564 3.64105 3.636 ;
		END
	END P19
	PIN P20
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 3.56895 3.564 3.64105 3.636 ;
		END
	END P20
	PIN P21
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 3.56895 3.564 3.64105 3.636 ;
		END
	END P21
	PIN P22
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 3.56895 3.564 3.64105 3.636 ;
		END
	END P22
	PIN P23
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 3.56895 3.564 3.64105 3.636 ;
		END
	END P23
	PIN P24
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 3.56895 3.564 3.64105 3.636 ;
		END
	END P24
	PIN P25
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 3.56895 3.564 3.64105 3.636 ;
		END
	END P25
	PIN P26
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 3.56895 3.564 3.64105 3.636 ;
		END
	END P26
	PIN P27
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 3.56895 3.564 3.64105 3.636 ;
		END
	END P27
	PIN P28
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 3.56895 3.564 3.64105 3.636 ;
		END
	END P28
	PIN P29
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 3.56895 3.564 3.64105 3.636 ;
		END
	END P29
	PIN P30
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 3.56895 3.564 3.64105 3.636 ;
		END
	END P30
	PIN P31
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 3.56895 3.564 3.64105 3.636 ;
		END
	END P31
	PIN P32
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 3.56895 3.564 3.64105 3.636 ;
		END
	END P32
	PIN P33
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 3.56895 3.564 3.64105 3.636 ;
		END
	END P33
	PIN P34
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 3.56895 3.564 3.64105 3.636 ;
		END
	END P34
	PIN P35
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 3.56895 3.564 3.64105 3.636 ;
		END
	END P35
	PIN P36
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 3.56895 3.564 3.64105 3.636 ;
		END
	END P36
	PIN P37
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 3.56895 3.564 3.64105 3.636 ;
		END
	END P37
	PIN P38
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 3.56895 3.564 3.64105 3.636 ;
		END
	END P38
	PIN P39
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 3.56895 3.564 3.64105 3.636 ;
		END
	END P39
	PIN P40
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 3.56895 3.564 3.64105 3.636 ;
		END
	END P40
	PIN P41
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 3.56895 3.564 3.64105 3.636 ;
		END
	END P41
	PIN P42
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 3.56895 3.564 3.64105 3.636 ;
		END
	END P42
	PIN P43
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 3.56895 3.564 3.64105 3.636 ;
		END
	END P43
	PIN P44
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 3.56895 3.564 3.64105 3.636 ;
		END
	END P44
	PIN P45
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 3.56895 3.564 3.64105 3.636 ;
		END
	END P45
	PIN P46
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 3.56895 3.564 3.64105 3.636 ;
		END
	END P46
	PIN P47
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 3.56895 3.564 3.64105 3.636 ;
		END
	END P47
	PIN P48
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 3.56895 3.564 3.64105 3.636 ;
		END
	END P48
	PIN P49
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 3.56895 3.564 3.64105 3.636 ;
		END
	END P49
	PIN P50
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 3.56895 3.564 3.64105 3.636 ;
		END
	END P50
	PIN P51
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 3.56895 3.564 3.64105 3.636 ;
		END
	END P51
	PIN P52
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 3.56895 3.564 3.64105 3.636 ;
		END
	END P52
	PIN P53
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 3.56895 3.564 3.64105 3.636 ;
		END
	END P53
END MAS68

MACRO MAS69
	CLASS CORE ;
	SIZE 9.85 BY 9.76 ;
	ORIGIN 0 0 ;
	SYMMETRY X ;
	SITE core 0 0 N DO 1 BY 1 STEP 0 0 ;
	PIN P1
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 4.87575 4.8312 4.97425 4.9288 ;
		END
	END P1
	PIN P2
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 4.87575 4.8312 4.97425 4.9288 ;
		END
	END P2
	PIN P3
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 4.87575 4.8312 4.97425 4.9288 ;
		END
	END P3
	PIN P4
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 4.87575 4.8312 4.97425 4.9288 ;
		END
	END P4
	PIN P5
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 4.87575 4.8312 4.97425 4.9288 ;
		END
	END P5
	PIN P6
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 4.87575 4.8312 4.97425 4.9288 ;
		END
	END P6
	PIN P7
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 4.87575 4.8312 4.97425 4.9288 ;
		END
	END P7
	PIN P8
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 4.87575 4.8312 4.97425 4.9288 ;
		END
	END P8
	PIN P9
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 4.87575 4.8312 4.97425 4.9288 ;
		END
	END P9
	PIN P10
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 4.87575 4.8312 4.97425 4.9288 ;
		END
	END P10
	PIN P11
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 4.87575 4.8312 4.97425 4.9288 ;
		END
	END P11
	PIN P12
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 4.87575 4.8312 4.97425 4.9288 ;
		END
	END P12
	PIN P13
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 4.87575 4.8312 4.97425 4.9288 ;
		END
	END P13
	PIN P14
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 4.87575 4.8312 4.97425 4.9288 ;
		END
	END P14
	PIN P15
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 4.87575 4.8312 4.97425 4.9288 ;
		END
	END P15
	PIN P16
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 4.87575 4.8312 4.97425 4.9288 ;
		END
	END P16
	PIN P17
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 4.87575 4.8312 4.97425 4.9288 ;
		END
	END P17
	PIN P18
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 4.87575 4.8312 4.97425 4.9288 ;
		END
	END P18
	PIN P19
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 4.87575 4.8312 4.97425 4.9288 ;
		END
	END P19
	PIN P20
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 4.87575 4.8312 4.97425 4.9288 ;
		END
	END P20
	PIN P21
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 4.87575 4.8312 4.97425 4.9288 ;
		END
	END P21
	PIN P22
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 4.87575 4.8312 4.97425 4.9288 ;
		END
	END P22
	PIN P23
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 4.87575 4.8312 4.97425 4.9288 ;
		END
	END P23
	PIN P24
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 4.87575 4.8312 4.97425 4.9288 ;
		END
	END P24
	PIN P25
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 4.87575 4.8312 4.97425 4.9288 ;
		END
	END P25
	PIN P26
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 4.87575 4.8312 4.97425 4.9288 ;
		END
	END P26
	PIN P27
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 4.87575 4.8312 4.97425 4.9288 ;
		END
	END P27
	PIN P28
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 4.87575 4.8312 4.97425 4.9288 ;
		END
	END P28
	PIN P29
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 4.87575 4.8312 4.97425 4.9288 ;
		END
	END P29
	PIN P30
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 4.87575 4.8312 4.97425 4.9288 ;
		END
	END P30
	PIN P31
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 4.87575 4.8312 4.97425 4.9288 ;
		END
	END P31
	PIN P32
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 4.87575 4.8312 4.97425 4.9288 ;
		END
	END P32
	PIN P33
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 4.87575 4.8312 4.97425 4.9288 ;
		END
	END P33
	PIN P34
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 4.87575 4.8312 4.97425 4.9288 ;
		END
	END P34
	PIN P35
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 4.87575 4.8312 4.97425 4.9288 ;
		END
	END P35
	PIN P36
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 4.87575 4.8312 4.97425 4.9288 ;
		END
	END P36
	PIN P37
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 4.87575 4.8312 4.97425 4.9288 ;
		END
	END P37
	PIN P38
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 4.87575 4.8312 4.97425 4.9288 ;
		END
	END P38
	PIN P39
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 4.87575 4.8312 4.97425 4.9288 ;
		END
	END P39
	PIN P40
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 4.87575 4.8312 4.97425 4.9288 ;
		END
	END P40
	PIN P41
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 4.87575 4.8312 4.97425 4.9288 ;
		END
	END P41
	PIN P42
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 4.87575 4.8312 4.97425 4.9288 ;
		END
	END P42
	PIN P43
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 4.87575 4.8312 4.97425 4.9288 ;
		END
	END P43
	PIN P44
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 4.87575 4.8312 4.97425 4.9288 ;
		END
	END P44
	PIN P45
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 4.87575 4.8312 4.97425 4.9288 ;
		END
	END P45
	PIN P46
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 4.87575 4.8312 4.97425 4.9288 ;
		END
	END P46
	PIN P47
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 4.87575 4.8312 4.97425 4.9288 ;
		END
	END P47
	PIN P48
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 4.87575 4.8312 4.97425 4.9288 ;
		END
	END P48
	PIN P49
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 4.87575 4.8312 4.97425 4.9288 ;
		END
	END P49
	PIN P50
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 4.87575 4.8312 4.97425 4.9288 ;
		END
	END P50
	PIN P51
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 4.87575 4.8312 4.97425 4.9288 ;
		END
	END P51
	PIN P52
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 4.87575 4.8312 4.97425 4.9288 ;
		END
	END P52
	PIN P53
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 4.87575 4.8312 4.97425 4.9288 ;
		END
	END P53
	PIN P54
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 4.87575 4.8312 4.97425 4.9288 ;
		END
	END P54
	PIN P55
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 4.87575 4.8312 4.97425 4.9288 ;
		END
	END P55
	PIN P56
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 4.87575 4.8312 4.97425 4.9288 ;
		END
	END P56
	PIN P57
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 4.87575 4.8312 4.97425 4.9288 ;
		END
	END P57
	PIN P58
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 4.87575 4.8312 4.97425 4.9288 ;
		END
	END P58
	PIN P59
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 4.87575 4.8312 4.97425 4.9288 ;
		END
	END P59
	PIN P60
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 4.87575 4.8312 4.97425 4.9288 ;
		END
	END P60
	PIN P61
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 4.87575 4.8312 4.97425 4.9288 ;
		END
	END P61
	PIN P62
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 4.87575 4.8312 4.97425 4.9288 ;
		END
	END P62
	PIN P63
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 4.87575 4.8312 4.97425 4.9288 ;
		END
	END P63
	PIN P64
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 4.87575 4.8312 4.97425 4.9288 ;
		END
	END P64
	PIN P65
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 4.87575 4.8312 4.97425 4.9288 ;
		END
	END P65
	PIN P66
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 4.87575 4.8312 4.97425 4.9288 ;
		END
	END P66
	PIN P67
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 4.87575 4.8312 4.97425 4.9288 ;
		END
	END P67
	PIN P68
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 4.87575 4.8312 4.97425 4.9288 ;
		END
	END P68
	PIN P69
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER metal1 ;
				RECT 4.87575 4.8312 4.97425 4.9288 ;
		END
	END P69
END MAS69

END LIBRARY

